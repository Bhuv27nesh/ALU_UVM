`define DATA_WIDTH 8
`define CMD_WIDTH 4

`define num_txns 2

`define SHIFT_WIDTH  $clog2(`DATA_WIDTH)
